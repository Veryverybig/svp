module mem(
    cpu_mem.tx cpu_mem
);

endmodule