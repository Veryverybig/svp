module cpu(
    cpu_mem.tx cpu_mem
);


endmodule